module gw_gao(
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[15] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[14] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[13] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[12] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[11] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[10] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[9] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[8] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[7] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[6] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[5] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[4] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[3] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[2] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[1] ,
    \pwm_top_dut/u_pwm_core_1/psc_preload_w[0] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[15] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[14] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[13] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[12] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[11] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[10] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[9] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[8] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[7] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[6] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[5] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[4] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[3] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[2] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[1] ,
    \pwm_top_dut/u_pwm_core_1/arr_preload_w[0] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[15] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[14] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[13] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[12] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[11] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[10] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[9] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[8] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[7] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[6] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[5] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[4] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[3] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[2] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[1] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[0] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[15] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[14] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[13] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[12] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[11] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[10] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[9] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[8] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[7] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[6] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[5] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[4] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[3] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[2] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[1] ,
    \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[0] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[15] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[14] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[13] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[12] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[11] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[10] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[9] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[8] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[7] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[6] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[5] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[4] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[3] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[2] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[1] ,
    \pwm_top_dut/u_pwm_core_1/cnt_val_w[0] ,
    \pwm_top_dut/u_pwm_core_1/cnt_en_w ,
    \pwm_top_dut/u_pwm_core_1/clk_psc_i ,
    \pwm_top_dut/u_pwm_core_1/ck_cnt_w ,
    \pwm_top_dut/u_pwm_core_1/pwm_ch1_a_o ,
    \pwm_top_dut/u_pwm_core_1/cnt_eq_cmp_ch1_start_w ,
    \pwm_top_dut/u_pwm_core_1/cnt_gt_cmp_ch1_start_w ,
    \pwm_top_dut/sys_soft_rst_i ,
    \pwm_top_dut/sys_hard_rst_i ,
    \pwm_top_dut/rst_n_i ,
    capture,
    clk_pwm,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \pwm_top_dut/u_pwm_core_1/psc_preload_w[15] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[14] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[13] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[12] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[11] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[10] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[9] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[8] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[7] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[6] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[5] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[4] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[3] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[2] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[1] ;
input \pwm_top_dut/u_pwm_core_1/psc_preload_w[0] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[15] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[14] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[13] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[12] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[11] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[10] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[9] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[8] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[7] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[6] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[5] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[4] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[3] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[2] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[1] ;
input \pwm_top_dut/u_pwm_core_1/arr_preload_w[0] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[15] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[14] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[13] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[12] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[11] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[10] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[9] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[8] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[7] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[6] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[5] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[4] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[3] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[2] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[1] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[0] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[15] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[14] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[13] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[12] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[11] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[10] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[9] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[8] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[7] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[6] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[5] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[4] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[3] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[2] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[1] ;
input \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[0] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[15] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[14] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[13] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[12] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[11] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[10] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[9] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[8] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[7] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[6] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[5] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[4] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[3] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[2] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[1] ;
input \pwm_top_dut/u_pwm_core_1/cnt_val_w[0] ;
input \pwm_top_dut/u_pwm_core_1/cnt_en_w ;
input \pwm_top_dut/u_pwm_core_1/clk_psc_i ;
input \pwm_top_dut/u_pwm_core_1/ck_cnt_w ;
input \pwm_top_dut/u_pwm_core_1/pwm_ch1_a_o ;
input \pwm_top_dut/u_pwm_core_1/cnt_eq_cmp_ch1_start_w ;
input \pwm_top_dut/u_pwm_core_1/cnt_gt_cmp_ch1_start_w ;
input \pwm_top_dut/sys_soft_rst_i ;
input \pwm_top_dut/sys_hard_rst_i ;
input \pwm_top_dut/rst_n_i ;
input capture;
input clk_pwm;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[15] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[14] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[13] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[12] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[11] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[10] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[9] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[8] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[7] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[6] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[5] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[4] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[3] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[2] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[1] ;
wire \pwm_top_dut/u_pwm_core_1/psc_preload_w[0] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[15] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[14] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[13] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[12] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[11] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[10] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[9] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[8] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[7] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[6] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[5] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[4] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[3] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[2] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[1] ;
wire \pwm_top_dut/u_pwm_core_1/arr_preload_w[0] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[15] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[14] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[13] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[12] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[11] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[10] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[9] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[8] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[7] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[6] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[5] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[4] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[3] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[2] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[1] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[0] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[15] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[14] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[13] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[12] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[11] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[10] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[9] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[8] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[7] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[6] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[5] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[4] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[3] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[2] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[1] ;
wire \pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[0] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[15] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[14] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[13] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[12] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[11] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[10] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[9] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[8] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[7] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[6] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[5] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[4] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[3] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[2] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[1] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_val_w[0] ;
wire \pwm_top_dut/u_pwm_core_1/cnt_en_w ;
wire \pwm_top_dut/u_pwm_core_1/clk_psc_i ;
wire \pwm_top_dut/u_pwm_core_1/ck_cnt_w ;
wire \pwm_top_dut/u_pwm_core_1/pwm_ch1_a_o ;
wire \pwm_top_dut/u_pwm_core_1/cnt_eq_cmp_ch1_start_w ;
wire \pwm_top_dut/u_pwm_core_1/cnt_gt_cmp_ch1_start_w ;
wire \pwm_top_dut/sys_soft_rst_i ;
wire \pwm_top_dut/sys_hard_rst_i ;
wire \pwm_top_dut/rst_n_i ;
wire capture;
wire clk_pwm;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i(capture),
    .trig1_i(\pwm_top_dut/sys_soft_rst_i ),
    .data_i({\pwm_top_dut/u_pwm_core_1/psc_preload_w[15] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[14] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[13] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[12] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[11] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[10] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[9] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[8] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[7] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[6] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[5] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[4] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[3] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[2] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[1] ,\pwm_top_dut/u_pwm_core_1/psc_preload_w[0] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[15] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[14] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[13] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[12] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[11] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[10] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[9] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[8] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[7] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[6] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[5] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[4] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[3] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[2] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[1] ,\pwm_top_dut/u_pwm_core_1/arr_preload_w[0] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[15] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[14] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[13] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[12] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[11] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[10] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[9] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[8] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[7] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[6] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[5] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[4] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[3] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[2] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[1] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_start_w[0] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[15] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[14] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[13] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[12] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[11] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[10] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[9] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[8] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[7] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[6] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[5] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[4] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[3] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[2] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[1] ,\pwm_top_dut/u_pwm_core_1/cmp_ch1_end_w[0] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[15] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[14] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[13] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[12] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[11] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[10] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[9] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[8] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[7] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[6] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[5] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[4] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[3] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[2] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[1] ,\pwm_top_dut/u_pwm_core_1/cnt_val_w[0] ,\pwm_top_dut/u_pwm_core_1/cnt_en_w ,\pwm_top_dut/u_pwm_core_1/clk_psc_i ,\pwm_top_dut/u_pwm_core_1/ck_cnt_w ,\pwm_top_dut/u_pwm_core_1/pwm_ch1_a_o ,\pwm_top_dut/u_pwm_core_1/cnt_eq_cmp_ch1_start_w ,\pwm_top_dut/u_pwm_core_1/cnt_gt_cmp_ch1_start_w ,\pwm_top_dut/sys_soft_rst_i ,\pwm_top_dut/sys_hard_rst_i ,\pwm_top_dut/rst_n_i }),
    .clk_i(clk_pwm)
);

endmodule
